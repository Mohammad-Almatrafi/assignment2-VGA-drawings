module tb_circles_datapath;



endmodule
