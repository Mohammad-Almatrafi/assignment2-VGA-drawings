
module tb_fillTheSreen_FSM;



endmodule
