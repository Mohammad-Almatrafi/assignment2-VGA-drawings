module tb_circles_controller;


endmodule
