
module tb_fillTheSreen_controller;



endmodule
