module tb_fillTheSreen_datapath;



endmodule
